
/*
 * Interfaces the camera to the rest of the system. Collects VGA frames from camera and writes it to the 2-PORT RAM block.
 * Documentation for all related to the camera (timing, configurations) can be found in the doc directory at the root of this repository	
 *
 *	Written by Ryan Song
 */
 
 module ov7670_driver();
 
 
 endmodule 
 
 
 /* Writes the data from the ov7670 camera to the 2-PORT RAM block */
 module ov7670_mem_ctrl();
	
 
 endmodule 