/*
 * This is the top level block for the embedded-cv project. 
 */
 
 module embedded_cv(  );
		
		
		
 
 endmodule 